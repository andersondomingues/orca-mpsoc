keep.me
