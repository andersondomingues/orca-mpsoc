fifo here
